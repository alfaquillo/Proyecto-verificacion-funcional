`timescale 1ns / 1ps

// =============================================================================
// Module: Template
// =============================================================================
// Descripción: Este modulo es una plantilla de formato 
//   
//
// Entradas:
//   
// Salidas:
//   
// Parámetros:
//   
// =============================================================================

module Template(

    );
endmodule
