`timescale 1ns / 1ps

// =============================================================================
// Module: 
// =============================================================================
// Descripción:
//   
//
// Entradas:
//   
//   
//   
//   
//
// Salidas:
//   
//
// Parámetros:
//   
//
// =============================================================================

module DecodificadorWR(WR, SEL, WE);

    input WR;
    input [3:0] SEL;
    output reg [11:0] WE;

    always @(*) 
    begin
        case ({WR, SEL})
            5'b10000: WE = 12'b000000000001;
            5'b10001: WE = 12'b000000000010;
            5'b10010: WE = 12'b000000000100;
            5'b10011: WE = 12'b000000001000;
            5'b10100: WE = 12'b000000010000;
            5'b10101: WE = 12'b000000100000;
            5'b10110: WE = 12'b000001000000;
            5'b10111: WE = 12'b000010000000;
            5'b11000: WE = 12'b000100000000;
            5'b11001: WE = 12'b001000000000;
            5'b11010: WE = 12'b010000000000;
            5'b11011: WE = 12'b100000000000;
            default:  WE = 12'b000000000000;
        endcase
    end

endmodule
