module Multiplexor6a1de16bits (A, B, C, D, E, F, SEL, OUT);

    input [15:0] A, B, C, D, E, F;
    input [2:0] SEL;
    output wire [15:0] OUT;

    assign OUT = (SEL == 3'd0) ? A :
                (SEL == 3'd1) ? B :
                (SEL == 3'd2) ? C :
                (SEL == 3'd3) ? D :
                (SEL == 3'd4) ? E :
                (SEL == 3'd5) ? F :
                16'd0;

endmodule